-------------------------------------------------------------------------------
-- Design: ALU / Entity / Project                                            --
--                                                                           --
-- Author : Sebastian Dichler                                                --
-- Date : 17. November 2017                                                  --
-- File : alu_entity.vhd                                                     --
-------------------------------------------------------------------------------


