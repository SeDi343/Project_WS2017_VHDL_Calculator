-------------------------------------------------------------------------------
-- Design: Testbench ALU / Project                                           --
--                                                                           --
-- Author : Sebastian Dichler                                                --
-- Date : 17. November 2017                                                  --
-- File : tb_alu.vhd                                                         --
-------------------------------------------------------------------------------


