-------------------------------------------------------------------------------
-- Design: CALC-CTRL / Entity / Project                                      --
--                                                                           --
-- Author : Sebastian Dichler                                                --
-- Date : 17. November 2017                                                  --
-- File : calc_entity_ctrl.vhd                                               --
-------------------------------------------------------------------------------


