-------------------------------------------------------------------------------
-- Design: Testbench CALC-CTRL / Project                                     --
--                                                                           --
-- Author : Sebastian Dichler                                                --
-- Date : 17. November 2017                                                  --
-- File : tb_calc_ctrl.vhd                                                   --
-------------------------------------------------------------------------------


