-------------------------------------------------------------------------------
-- Design: Testbench IO-CTRL / Project                                       --
--                                                                           --
-- Author : Sebastian Dichler                                                --
-- Date : 17. November 2017                                                  --
-- File : tb_io_ctrl.vhd                                                     --
-------------------------------------------------------------------------------


